module sequencer(clk, flag, out);
parameter N=2;

endmodule