module sequencer_test(clk, led);
input clk;
output [] led;
endmodule